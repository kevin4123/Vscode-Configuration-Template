/* @wavedrom counter waveform
{
  signal: [
    { name: "clk",   wave: "p.p.p.p.p.p.p.p" },
    { name: "rst",   wave: "10..........." },
    { name: "count", wave: "x============", data: ["0", "1", "2", "3", "4", "5", "6","7","8","9","10","11"] }
  ],
  head: {
    text: "4-bit Counter Waveform",
    tick: 0,
  },
  foot: {
    text: "Counter counts on each positive clock edge when reset is low",
    tick: 0,
  }
}
*/

module counter (
    input  wire clk,
    input  wire rst,
    output reg [3:0] count
);

    always @(posedge clk or posedge rst) begin
        if (rst)
            count <= 4'b0000;
        else
            count <= count + 1;
    end
endmodule
